module control_logic #() (); 
endmodule
