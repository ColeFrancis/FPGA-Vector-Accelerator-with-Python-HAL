module top #() ();
endmodule
